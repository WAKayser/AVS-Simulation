module fsmTb;

reg clock, reset;
reg signed serial;
wire eventDetected;

topLevel topLevel (.clock(clock),.reset(reset),.serial(serial),.eventDetected(eventDetected),.uart_out(uart_out));

initial begin
	clock = 0;
	reset = 1;
	serial = 0;

	#100 reset = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;
	#10000 serial = 1;
	#1000 serial = 0;



end

always
#5 clock =! clock;


endmodule